----------------------------------------------------------------------------------
-- Project Name: Frecuency Counter 
-- Target Devices: Spartan 3
-- Engineers: �ngel Larra�aga Muro
-- 			 Nicol�s Jurado Jim�nez
-- 			 Gonzalo Matarrubia Gonzalez
-- License: All files included in this proyect are licensed under a Creative Commons Attribution-ShareAlike 4.0 International License 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
 
entity clk_mod is
    Port (
        entrada: in  STD_LOGIC;
        reset  : in  STD_LOGIC;
        salida : out STD_LOGIC
    );
end clk_mod;
 
architecture Behavioral of clk_mod is
    signal temporal: STD_LOGIC;
    signal contador: integer range 0 to 150000 := 0;
begin
    divisor_frecuencia: process (reset, entrada) begin
        if (reset = '1') then
            temporal <= '0';
            contador <= 0;
        elsif rising_edge(entrada) then
            if (contador = 25000) then 			--ESTA VARIABLE ES LA QUE HACE QUE SE MODIFICA LA FRECUENCIA. HAY QUE DIVIDIR LA DEL RELOJ DE LA TARJETA ENTRE LA DESEADA Y DIVIDIRLA ENTRE 2 (semiperiodo).
                temporal <= NOT(temporal);
                contador <= 0;
            else
                contador <= contador+1;
            end if;
        end if;
    end process;
     
    salida <= temporal;
end Behavioral;